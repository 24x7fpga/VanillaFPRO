kiran@SuperComp.1334:1716351544